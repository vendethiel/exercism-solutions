module main

fn hello() string {
	return 'Hello, World!'
}
